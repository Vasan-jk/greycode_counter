/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none
/*
module tt_um_example (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // All output pins must be assigned. If not used, assign to 0.
  assign uo_out  = ui_in + uio_in;  // Example: ou_out is the sum of ui_in and uio_in
  assign uio_out = 0;
  assign uio_oe  = 0;

  // List all unused inputs to prevent warnings
  wire _unused = &{ena, clk, rst_n, 1'b0};

endmodule
*/

// gray_counter.v
// Fixed 8-bit Gray Code Counter
/*
module gray_counter (
    input  wire       clk,    // clock
    input  wire       rst_n,  // active-low reset
    output reg [7:0]  gray    // Gray code output
);

    reg [7:0] binary;  // internal binary counter

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            binary <= 8'd0;
            gray   <= 8'd0;
        end else begin
            binary <= binary + 1'b1;          // increment binary counter
            gray   <= binary ^ (binary >> 1); // convert to Gray code
        end
    end

endmodule
*/
// 8-bit Gray Code Counter for TinyTapeout
module tt_um_gray_counter (
    input  wire [7:0] ui_in,    // unused user inputs
    output wire [7:0] uo_out,   // Gray code output
    input  wire [7:0] uio_in,   // unused bidirectional inputs
    output wire [7:0] uio_out,  // unused bidirectional outputs
    output wire [7:0] uio_oe,   // unused output enables
    input  wire       clk,      // global clock
    input  wire       rst_n     // global reset (active low)
);

    reg [7:0] binary;
    reg [7:0] gray;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            binary <= 8'b0;
            gray   <= 8'b0;
        end else begin
            binary <= binary + 1'b1;
            gray   <= binary ^ (binary >> 1);
        end
    end

    // Drive outputs
    assign uo_out  = gray;

    // Not using bidirectional IOs
    assign uio_out = 8'b0;
    assign uio_oe  = 8'b0;

endmodule

